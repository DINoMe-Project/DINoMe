module NBDTLB( // @[:example.TestHarness.TinyBoomConfig1.fir@214641.2]
  input         clock, // @[:example.TestHarness.TinyBoomConfig1.fir@214642.4]
  input         reset, // @[:example.TestHarness.TinyBoomConfig1.fir@214643.4]
  output        io_req_0_ready, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_req_0_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_req_0_bits_vaddr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_req_0_bits_passthrough, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_req_0_bits_size, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [4:0]  io_req_0_bits_cmd, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_miss_rdy, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_miss, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output [31:0] io_resp_0_paddr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_pf_ld, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_pf_st, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_ae_ld, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_ae_st, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_ma_ld, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_ma_st, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_resp_0_cacheable, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_sfence_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_sfence_bits_rs1, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_sfence_bits_rs2, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_sfence_bits_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_req_ready, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_ptw_req_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output        io_ptw_req_bits_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_ae, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_d, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_g, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_u, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_pte_v, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_level, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_resp_bits_homogeneous, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_ptbr_mode, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_status_dprv, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_status_mxr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_status_sum, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_0_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_0_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_0_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_0_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_1_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_1_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_1_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_1_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_2_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_2_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_2_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_2_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_3_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_3_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_3_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_3_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_4_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_4_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_4_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_4_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_5_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_5_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_5_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_5_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_6_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_6_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_6_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_6_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_7_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_7_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_7_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_ptw_pmp_7_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input  [31:0] io_ptw_pmp_7_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
  input         io_kill // @[:example.TestHarness.TinyBoomConfig1.fir@214644.4]
);
assign io_resp_0_paddr=io_req_0_bits_vaddr;
assign io_req_0_ready = io_req_0_valid;
assign io_resp_0_miss= ~io_req_0_valid;
assign io_miss_rdy =1'b0;
assign io_resp_0_cacheable=1'b1;
assign io_resp_0_ae_st=1'b0;
assign io_resp_0_ae_ld=1'b0;
assign io_resp_0_ma_st=1'b0;
assign io_resp_0_ma_ld=1'b0;
assign io_resp_0_pf_ld=1'b0;
assign io_resp_0_pf_st=1'b0;
assign io_ptw_req_valid=1'b0;
assign io_ptw_req_bits_bits_valid=1'b0;
assign io_ptw_req_bits_bits_addr=io_req_0_bits_vaddr[31:12];
endmodule
module TLB( // @[:example.TestHarness.TinyBoomConfig1.fir@146269.2]
  input         clock, // @[:example.TestHarness.TinyBoomConfig1.fir@146270.4]
  input         reset, // @[:example.TestHarness.TinyBoomConfig1.fir@146271.4]
  output        io_req_ready, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_req_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_req_bits_vaddr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output        io_resp_miss, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output [31:0] io_resp_paddr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output        io_resp_pf_inst, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output        io_resp_ae_inst, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output        io_resp_cacheable, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_sfence_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_sfence_bits_rs1, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_sfence_bits_rs2, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_sfence_bits_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_req_ready, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output        io_ptw_req_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_valid, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_ae, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_d, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_g, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_u, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_pte_v, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_level, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_resp_bits_homogeneous, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_ptbr_mode, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_status_prv, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_0_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_0_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_0_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_0_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_1_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_1_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_1_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_1_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_2_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_2_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_2_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_2_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_3_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_3_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_3_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_3_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_4_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_4_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_4_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_4_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_5_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_5_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_5_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_5_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_6_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_6_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_6_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_6_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_7_cfg_l, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_7_cfg_x, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_7_cfg_w, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input         io_ptw_pmp_7_cfg_r, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
  input  [31:0] io_ptw_pmp_7_mask // @[:example.TestHarness.TinyBoomConfig1.fir@146272.4]
);

assign io_req_ready = io_req_valid;
assign io_resp_miss = ~io_req_valid;
assign io_resp_paddr=io_req_bits_vaddr;
assign io_resp_pf_inst=1'h0;
assign io_resp_ae_inst=1'h0;
assign io_resp_cacheable=1'b1;
assign io_ptw_req_valid=1'b0;
assign io_ptw_req_bits_bits_addr=io_req_bits_vaddr[31:12];
endmodule

module TLB_new( // @[:example.TestHarness.TinyBoomConfig8.fir@65045.2]
  input         clock, // @[:example.TestHarness.TinyBoomConfig8.fir@65046.4]
  input         reset, // @[:example.TestHarness.TinyBoomConfig8.fir@65047.4]
  output        io_req_ready, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_req_valid, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_req_bits_vaddr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output        io_resp_miss, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output [31:0] io_resp_paddr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output        io_resp_pf_inst, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output        io_resp_ae_inst, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output        io_resp_cacheable, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_sfence_valid, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_sfence_bits_rs1, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_sfence_bits_rs2, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_sfence_bits_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_req_ready, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output        io_ptw_req_valid, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  output [19:0] io_ptw_req_bits_bits_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_valid, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_ae, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [53:0] io_ptw_resp_bits_pte_ppn, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_d, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_g, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_u, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_pte_v, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_level, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_resp_bits_homogeneous, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_ptbr_mode, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_status_prv, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_0_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_0_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_0_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_0_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_0_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_0_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_0_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_1_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_1_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_1_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_1_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_1_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_1_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_1_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_2_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_2_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_2_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_2_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_2_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_2_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_2_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_3_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_3_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_3_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_3_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_3_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_3_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_3_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_4_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_4_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_4_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_4_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_4_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_4_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_4_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_5_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_5_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_5_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_5_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_5_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_5_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_5_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_6_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_6_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_6_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_6_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_6_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_6_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_6_mask, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_7_cfg_l, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [1:0]  io_ptw_pmp_7_cfg_a, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_7_cfg_x, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_7_cfg_w, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input         io_ptw_pmp_7_cfg_r, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [29:0] io_ptw_pmp_7_addr, // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
  input  [31:0] io_ptw_pmp_7_mask // @[:example.TestHarness.TinyBoomConfig8.fir@65048.4]
);
assign io_req_ready = io_req_valid;
assign io_resp_miss = ~io_req_valid;
assign io_resp_paddr=io_req_bits_vaddr;
assign io_resp_pf_inst=1'h0;
assign io_resp_ae_inst=1'h0;
assign io_resp_cacheable=1'b1;
assign io_ptw_req_valid=1'b0;
assign io_ptw_req_bits_bits_addr=io_req_bits_vaddr[31:12];
endmodule
